`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:48:35 11/11/2019 
// Design Name: 
// Module Name:    controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module controller(
    input [5:0] opc,
    input [5:0] func,
    output regdst,
    output alusrc,
    output memtoreg,
    output regwrite,
    output memwrite,
    output memread,
    output extop,
    output luiop,
    output [2:0] aluop,
    output [2:0] npc_slc,
    output jalop,
	 output jalrop,
	 output sraop
    );
	 wire addu,subu,ori,lw,sw,beq,lui,jal,jr;
	 
	 assign addu = ((opc==6'b000000)&&(func==6'b100001));
	 assign subu = ((opc==6'b000000)&&(func==6'b100011));
	 assign ori = (opc==6'b001101);
	 assign lw = (opc==6'b100011);
	 assign sw = (opc==6'b101011);
	 assign beq = (opc==6'b000100);
	 assign lui = (opc==6'b001111);
	 assign jal = (opc==6'b000011);
	 assign jr = ((opc==6'b000000)&&(func==6'b001000));
	 assign j = (opc==6'b000010);
	 assign jalr = ((opc==6'b000000)&&(func==6'b001001));
	 assign sra = ((opc==6'b000000)&&(func==6'b000011));
	 
	 assign regdst = addu || subu || sra;
	 assign alusrc = ori || lw || sw || lui;
	 assign memtoreg = lw;
	 assign regwrite = addu || jal || subu || lw || lui || ori || jalr || sra;
	 assign memwrite = sw;
	 assign memread = lw;
	 assign extop = sw || lw || beq;
	 assign luiop = lui;
	 assign jalop = jal;
	 assign jalrop = jalr;
	 assign sraop = sra;
	 
	 assign aluop[2] = 0;
	 assign aluop[1] = addu || subu || lw || sw || lui;
	 assign aluop[0] = subu || ori;
	 
	 assign npc_slc[2] = jr || jalr; 
	 assign npc_slc[1] = jal || j ;
	 assign npc_slc[0] = jal || beq || jalr;
	 

endmodule
